netcdf x2b_h2o_ion_v1 {
  // global attributes
  :name = "x2b_h2o_ion_v1<5>";
  :C6_XH =  5.681559999999999e+02; // kcal/mol * A^6
  :C6_XO =  1.294680000000000e+03; // kcal/mol * A^6
  :C8_XH =  0.000000000000000e+00; // kcal/mol * A^8
  :C8_XO =  0.000000000000000e+00; // kcal/mol * A^8
  :d6_XH =  2.930890000000000e+00; // A^(-1)
  :d6_XO =  2.719380000000000e+00; // A^(-1)
  :d8_XH =  2.000000000000000e+00; // A^(-1)
  :d8_XO =  2.000000000000000e+00; // A^(-1)
  :k_HH_intra =  7.952670334647889e-01; // A^(-1)
  :k_OH_intra =  3.669544414655080e-01; // A^(-1)
  :k_XH_coul =  2.836253042727388e-01; // A^(-1)
  :k_XO_coul =  3.693558640786222e-01; // A^(-1)
  :k_xlp_main =  3.687700750039854e-01; // A^(-1)
  :d_HH_intra =  1.999999814890842e+00; // A^(-1)
  :d_OH_intra =  1.309170470030335e+00; // A^(-1)
  :d_XH_coul =  5.914094693840913e+00; // A^(-1)
  :d_XO_coul =  6.941993233395817e+00; // A^(-1)
  :d_xlp_main =  5.557092273485791e+00; // A^(-1)
  :in_plane_gamma =  3.762643956966366e-03;
  :out_of_plane_gamma =  9.221730898707543e-01;
  :r2i =  6.000000000000000e+00; // A
  :r2f =  7.000000000000000e+00; // A
  dimensions:
  poly = 429;
  variables:
    double poly(poly);
data:
poly =
 1.148769522971932e+02, // 0
-2.773230726991214e+02, // 1
 1.827078013468585e+01, // 2
 1.392387016304614e+02, // 3
-3.543937376542597e+02, // 4
-4.788932246721681e+01, // 5
 3.481270393056712e+02, // 6
-6.377371891853971e+02, // 7
-1.434213914638941e+02, // 8
-1.669483446893566e+01, // 9
-3.346122327292023e+02, // 10
-9.405921827092223e+00, // 11
-1.811425870210874e+02, // 12
-2.901047316502409e+02, // 13
-1.540200309952160e+02, // 14
-5.329377963408669e+01, // 15
-2.543637871643261e+01, // 16
 2.369450396732275e+02, // 17
 5.100420041747400e+02, // 18
 1.637358637520869e+02, // 19
 1.896175393139902e+02, // 20
-1.809182643635956e+02, // 21
-4.559721866561475e+01, // 22
 1.736985553316242e+02, // 23
 2.383489780642338e+02, // 24
 1.298843554056843e+02, // 25
 1.959466931005129e+02, // 26
-2.733371202853143e+01, // 27
-1.427079175611695e+01, // 28
-9.695294902699514e+00, // 29
-2.388203116803058e+02, // 30
-4.428511991508392e+01, // 31
 1.138115726037502e+02, // 32
 3.345609988242910e+01, // 33
 3.486326778990320e+02, // 34
 1.795611168334411e+01, // 35
-9.298896284954937e+01, // 36
-1.198736948163496e+01, // 37
 5.106356634337293e+01, // 38
-3.183411591578625e+02, // 39
 4.611685851864881e+01, // 40
 2.935757833512388e+02, // 41
-8.225562756834988e+01, // 42
-3.004280073051667e+02, // 43
 1.399028231126495e+02, // 44
-7.384308588145628e+01, // 45
 5.619597271486090e+01, // 46
 1.178389088868073e+03, // 47
-1.063226851316105e+02, // 48
 3.846787354466377e+02, // 49
 4.886571456843810e+01, // 50
-1.389924210899761e+02, // 51
-8.000272288343858e+00, // 52
-8.840846846371411e+00, // 53
 3.384116735813686e+02, // 54
 2.288646475592941e+02, // 55
-1.416969357419378e+02, // 56
-1.079211809836504e+01, // 57
-6.886951633066723e+00, // 58
-2.587880889121563e+02, // 59
 9.959730634903343e+01, // 60
 3.701308203675230e+01, // 61
 2.918291265575431e+01, // 62
 2.240033900886754e+02, // 63
 3.417831104637669e+01, // 64
 1.609368831363900e+02, // 65
 3.481728160027019e+02, // 66
 1.506067520281869e+01, // 67
-4.060287901080621e+01, // 68
 4.039634970432867e+01, // 69
-1.677142520167795e+01, // 70
-2.563091637785741e+01, // 71
 4.177221727382538e+02, // 72
-1.029233843619212e+02, // 73
 2.609061279287321e+02, // 74
 1.319184978370535e+02, // 75
-5.707005542736367e+01, // 76
-9.087282555351493e+00, // 77
-7.216428394853735e+02, // 78
 3.918397496833502e+01, // 79
 1.325220149204583e+02, // 80
-6.705334213482280e+01, // 81
 4.838027488738896e+01, // 82
 5.337675079110923e+01, // 83
 1.285067935868455e+01, // 84
 5.782081505373394e+01, // 85
 1.057169846084842e+01, // 86
 2.330629498219623e+01, // 87
-1.457184075610011e+02, // 88
 5.500266003389308e+01, // 89
-9.015220961283853e+01, // 90
-3.379570812520808e+02, // 91
-1.664017836343734e+02, // 92
 1.010267064832749e+01, // 93
 3.159432042901072e+02, // 94
 2.731384069552552e+00, // 95
-1.707535931830466e+01, // 96
 2.123432652862337e+01, // 97
 1.008565155326918e+02, // 98
 1.781493116943984e+02, // 99
-2.329441677621762e+02, // 100
-2.280388846745338e+01, // 101
-3.375072410101278e+01, // 102
 8.953594923964322e+01, // 103
-2.586840052853664e+01, // 104
-3.677873928569151e+02, // 105
 1.119123268293022e+01, // 106
-2.681676365620640e+01, // 107
 2.062966206262750e+01, // 108
 6.839486370960344e+02, // 109
-8.656616762047805e+01, // 110
 1.570578318100126e+01, // 111
-2.903434470445363e+02, // 112
-6.467586290635420e+01, // 113
-3.345669961313124e+02, // 114
-5.773108495138027e+00, // 115
 5.565647160788554e+00, // 116
-7.014078365103826e+01, // 117
-8.721229396247681e+01, // 118
-2.283364352213266e+02, // 119
-1.252041142827894e+01, // 120
-8.162446839448656e+01, // 121
 8.646998412935514e+01, // 122
 3.534885587499693e+00, // 123
-1.433203611752304e+01, // 124
 5.714893144903001e+00, // 125
 1.406875319524373e+01, // 126
-6.024747243022416e+01, // 127
-1.139102133817977e+01, // 128
-5.283478651529086e+01, // 129
 4.914450028329219e+01, // 130
 2.703500482104002e+01, // 131
-3.358141400035345e+01, // 132
-8.723168136019599e+02, // 133
 1.337726203635031e+02, // 134
 9.481344757477048e+01, // 135
 3.038708579275047e+01, // 136
 1.027816874091094e+03, // 137
-7.701909436455724e+02, // 138
-1.206731756029336e+02, // 139
-6.063798778298574e+00, // 140
 4.760623437982876e+01, // 141
 1.041485723698920e+01, // 142
 1.357884939436762e+02, // 143
 9.328926192113304e+00, // 144
-4.737647383608125e+01, // 145
-1.884061104801030e+02, // 146
-7.943057905924233e+01, // 147
 2.188953027249171e+02, // 148
 1.298078627915482e+02, // 149
-1.253961760422727e+02, // 150
 2.669007647967912e-01, // 151
 7.147033469439430e+01, // 152
 1.620314864022881e+02, // 153
 3.798774102490260e+00, // 154
 5.459705548251652e+01, // 155
-5.106099121505791e+02, // 156
-2.850620590777012e+01, // 157
-1.885978523416164e+02, // 158
 4.229823815329361e+01, // 159
 1.546564377044440e+02, // 160
-1.117156682655241e+02, // 161
-2.570166647031470e+02, // 162
-1.853191304224521e+02, // 163
-5.387050599225936e+01, // 164
 2.868766809850792e+02, // 165
-1.279324939946467e+02, // 166
-2.649231919344887e+02, // 167
-1.140401568224698e+02, // 168
-1.230599105479334e+02, // 169
-1.281524682620779e+02, // 170
-1.932777173932515e+01, // 171
 3.310965813859586e+02, // 172
-5.542895985264259e+02, // 173
-2.370209462461247e+01, // 174
-1.444521942656079e+02, // 175
-6.829870723785189e+01, // 176
-6.887199461676778e+01, // 177
 1.972881192395792e+02, // 178
-1.448108997519860e+02, // 179
 1.780133513151946e+02, // 180
-3.219191273740833e+02, // 181
-8.496263216416243e+01, // 182
 4.774279799015682e+01, // 183
 5.239999192094893e+01, // 184
 8.359481538763937e+01, // 185
-3.102057756434187e+00, // 186
 1.741948941202592e+02, // 187
-1.109748261916130e+02, // 188
 1.039221233261241e+01, // 189
-1.044819240934761e+02, // 190
 1.560755188881533e+01, // 191
-1.112545720413457e+02, // 192
-2.875830940812587e+01, // 193
-1.832402800118280e+02, // 194
 4.931212308940081e-01, // 195
 3.263696640970849e+00, // 196
 1.586791486114863e+02, // 197
 1.401309135420372e+02, // 198
-6.961550114291054e+00, // 199
 6.663133848315468e+00, // 200
 4.323263823387389e+01, // 201
-8.457720930279082e+00, // 202
 1.086059942152274e+01, // 203
-4.372390965886945e+00, // 204
-4.641207358943296e+01, // 205
 1.838575441249651e+01, // 206
-2.062846323839168e+01, // 207
-1.130946646149037e+01, // 208
 8.753879332220089e+01, // 209
 2.928276805231274e+01, // 210
 3.124304411105750e+01, // 211
-2.552317776578041e+01, // 212
 3.700575231702040e+01, // 213
-1.942279607219181e+01, // 214
 5.276925924213560e+00, // 215
 5.317471242562561e+01, // 216
 3.281111321828956e+02, // 217
-2.097146044480340e+01, // 218
-2.461602054118764e+01, // 219
 9.024790212526024e+01, // 220
-3.906503189218778e+01, // 221
-5.992682895020629e+01, // 222
-1.896388871297952e+01, // 223
-4.576152299348663e+00, // 224
-2.059488909670012e+01, // 225
 2.262688503327740e+01, // 226
-1.040503300826663e+01, // 227
 6.063274349299164e+01, // 228
-5.476540156533190e+00, // 229
-4.587224859937470e+01, // 230
 2.965449410156635e+02, // 231
 2.694826419763689e+01, // 232
-2.444340493144963e-01, // 233
 4.868577418071524e+00, // 234
 8.990402329935202e+00, // 235
 3.106022937891999e+02, // 236
-6.485667868589720e+00, // 237
 5.641371064387402e+00, // 238
-1.008045347254097e+01, // 239
-1.268207106746162e+01, // 240
 5.662372036810094e+01, // 241
 2.875084285145348e+01, // 242
-8.143941772364213e-01, // 243
-1.352864949406492e+01, // 244
-3.412984705403661e+01, // 245
 6.099970653155969e+00, // 246
 5.397198586546182e+01, // 247
 1.625144744038886e+01, // 248
 7.599976028679833e+00, // 249
-5.217166607294051e+01, // 250
 1.067236565008029e+00, // 251
-1.368872039087096e+01, // 252
-1.237032130024221e+02, // 253
-1.162686437889927e+01, // 254
-5.131970012324498e+00, // 255
 1.758603614235379e+02, // 256
 3.663384968441732e+01, // 257
-1.269734923169290e+01, // 258
 4.254380043484828e+01, // 259
 8.863976296754862e+00, // 260
 9.995614405441455e+01, // 261
 3.793527303867462e+01, // 262
-6.968119143717601e+00, // 263
-3.017916849165569e+01, // 264
-8.352303011778671e+00, // 265
 8.580288279937216e+00, // 266
-4.152630900138563e+01, // 267
-3.682000969235144e+01, // 268
-2.466045733896760e+01, // 269
-1.063043597934746e+02, // 270
-1.520203602213399e+01, // 271
-9.789796707495297e+00, // 272
 2.522417658762323e+01, // 273
-9.899569182663404e+00, // 274
-2.500778116830504e+01, // 275
 1.678409187239478e+01, // 276
-2.790005621282157e+01, // 277
 1.282594046519141e+02, // 278
-1.311711046109752e+01, // 279
-1.081477919012787e+01, // 280
-3.266610573530381e+01, // 281
 1.336527757778771e+01, // 282
-3.849178690423969e+00, // 283
 1.375097631424553e+01, // 284
 1.546472671136714e+00, // 285
 1.408489364545349e+02, // 286
-3.399167146512315e+01, // 287
 1.220584736924130e+02, // 288
 6.921909069514521e+01, // 289
-1.541854556397614e+01, // 290
-1.121683848519438e+01, // 291
-9.242430137881306e+01, // 292
 2.628408813066963e+00, // 293
-7.814789205760461e+01, // 294
 4.990575271723984e+00, // 295
 2.242325011070997e+01, // 296
-2.623474720305492e+02, // 297
 6.619640899108076e+00, // 298
-1.851266224027469e+01, // 299
 4.029454521727645e+01, // 300
-2.759983421798458e+00, // 301
-1.728167246766074e+00, // 302
-2.424292052728002e+02, // 303
-2.367667715221609e+01, // 304
-1.876198055462046e+02, // 305
-3.348194716549535e+00, // 306
 1.781243256485856e+01, // 307
 1.714765932860531e+02, // 308
 1.022496295069972e+01, // 309
 2.049319192106086e+02, // 310
-2.590315159006037e-01, // 311
-5.619827849628722e+01, // 312
-7.388918007227944e+01, // 313
-4.817616823928957e+00, // 314
 2.326785371460746e+00, // 315
 6.489031709802128e-01, // 316
 1.406158974433800e+01, // 317
-1.654667756391876e+00, // 318
 1.911775297265568e+01, // 319
-1.067786109390064e+02, // 320
 1.227641372085565e+01, // 321
 4.051469528739763e+00, // 322
-5.053892485705552e-01, // 323
 2.378888869936005e+01, // 324
-3.352250900843055e+01, // 325
-3.225766823141835e+01, // 326
-3.979634244415261e+01, // 327
-2.483585958374013e+01, // 328
-6.781421883778988e+00, // 329
 3.319870346003055e+01, // 330
 1.120586308603971e+02, // 331
-5.909233970862215e+00, // 332
 2.882230188200199e+01, // 333
 3.383547407485854e+01, // 334
-1.536743154204077e+01, // 335
 1.658523163566573e+01, // 336
-2.038831431215415e+01, // 337
 4.918959454655425e+01, // 338
 9.255618087520217e+01, // 339
 6.823492437749704e+00, // 340
-2.486279258926865e+00, // 341
 3.512070169200672e+01, // 342
 8.276298300902290e+01, // 343
 2.886948695746750e+00, // 344
-6.263508756304613e+01, // 345
 1.858070177354850e+01, // 346
 3.785461296096628e-01, // 347
 9.500823267075153e+01, // 348
 4.319414915742287e+00, // 349
 2.768879558267599e+01, // 350
-1.007141694321548e+01, // 351
 3.460815668996207e-01, // 352
-2.575480686473782e+01, // 353
 5.300716230333460e-01, // 354
 3.077891657909914e+02, // 355
 3.820408272122957e+01, // 356
 1.110648456196821e+01, // 357
 2.903639161993504e+02, // 358
-3.090515612059465e+00, // 359
 3.049170795430189e+02, // 360
-1.575710833651697e+00, // 361
-2.207182752692426e+01, // 362
-3.221504832613083e+01, // 363
 5.549706133232642e+01, // 364
 5.499564412381432e+00, // 365
-8.828859593923490e+00, // 366
-8.260904514927211e+01, // 367
 4.553657496482112e+01, // 368
 4.476021393925404e+01, // 369
-1.440628717503907e+00, // 370
-2.160596957012654e+01, // 371
 1.175446857335780e+02, // 372
 1.653861451581694e+00, // 373
 1.232700279138528e+01, // 374
 1.640760365353830e+02, // 375
 1.507624250051121e+01, // 376
-1.903561373928230e+01, // 377
 1.186475009234863e+01, // 378
 7.508451382944173e+00, // 379
-1.475904433573388e+01, // 380
 6.348715414739159e+01, // 381
 2.967420881611330e+01, // 382
 1.487294989194473e+01, // 383
-2.448899774129269e+01, // 384
 4.613419989482298e+01, // 385
 1.770314745535570e+00, // 386
-1.724754313934627e+02, // 387
 5.905479975172500e+01, // 388
 3.154443844135095e+01, // 389
-6.390132460405413e+02, // 390
-4.374391071346894e+02, // 391
 6.648263057930022e+01, // 392
-1.172060513462072e+00, // 393
-3.105607408856294e+01, // 394
-1.193486725173444e+01, // 395
-1.211627272133822e+02, // 396
-4.440307767540166e+00, // 397
 3.763693799360639e+00, // 398
-1.712025091780114e+02, // 399
 8.392696387372299e+00, // 400
 9.491484482160464e-01, // 401
-3.756131296714052e+00, // 402
 1.693948749381030e+01, // 403
 3.325063116325246e-01, // 404
 6.298214145684563e-01, // 405
 3.598871686954166e+01, // 406
 1.176906374533055e+01, // 407
-3.389957220576565e+02, // 408
-7.762765833362065e-01, // 409
-1.673005286087509e+00, // 410
-8.411998204489188e+01, // 411
-2.619653119920854e-01, // 412
 2.535155337193745e+01, // 413
 1.529482938535785e+01, // 414
-7.016189695203325e+00, // 415
-3.964555485076855e+01, // 416
 1.301629246558452e+00, // 417
 5.386131410693063e+02, // 418
-1.836567069804440e+01, // 419
 2.433060770970746e+00, // 420
-3.028635009467761e+02, // 421
 1.340981467914506e+01, // 422
-1.023930471155378e+01, // 423
 1.796950315414689e+01, // 424
 1.598791759505597e+01, // 425
-2.272672877280680e+00, // 426
-3.398291031027740e+01, // 427
 2.973014615468740e+01; // 428

}
